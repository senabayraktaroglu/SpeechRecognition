

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity hamming_rom is
--  Port ( );
port(clk: in std_logic;
    address: in integer range 0 to 511;
     data: out std_logic_vector(15 downto 0));
end hamming_rom;

architecture Behavioral of hamming_rom is
    type rom_array is array (0 to 511) of std_logic_vector (15 downto 0);
    constant rom: rom_array := (
    "0000000000001000",--1
    "0000000000001000",--2
    "0000000000001000",--3
    "0000000000001000",--4
    "0000000000001000",--5
    "0000000000001000",--6
    "0000000000001000",--7
    "0000000000001000",--8
    "0000000000001000",--9
    "0000000000001000",--10
    "0000000000001000",--11
    "0000000000001000",--12
    "0000000000001000",--13
    "0000000000001001",--14
    "0000000000001001",--15
    "0000000000001001",--16
    "0000000000001001",--17
    "0000000000001001",--18
    "0000000000001001",--19
    "0000000000001001",--20
    "0000000000001001",--21
    "0000000000001010",--22
    "0000000000001010",--23
    "0000000000001010",--24
    "0000000000001010",--25
    "0000000000001010",--26
    "0000000000001010",--27
    "0000000000001011",--28
    "0000000000001011",--29
    "0000000000001011",--30
    "0000000000001011",--31
    "0000000000001011",--32
    "0000000000001100",--33
    "0000000000001100",--34
    "0000000000001100",--35
    "0000000000001100",--36
    "0000000000001100",--37
    "0000000000001101",--38
    "0000000000001101",--39
    "0000000000001101",--40
    "0000000000001101",--41
    "0000000000001110",--42
    "0000000000001110",--43
    "0000000000001110",--44
    "0000000000001111",--45
    "0000000000001111",--46
    "0000000000001111",--47
    "0000000000001111",--48
    "0000000000010000",--49
    "0000000000010000",--50
    "0000000000010000",--51
    "0000000000010001",--52
    "0000000000010001",--53
    "0000000000010001",--54
    "0000000000010010",--55
    "0000000000010010",--56
    "0000000000010010",--57
    "0000000000010011",--58
    "0000000000010011",--59
    "0000000000010100",--60
    "0000000000010100",--61
    "0000000000010100",--62
    "0000000000010101",--63
    "0000000000010101",--64
    "0000000000010110",--65
    "0000000000010110",--66
    "0000000000010110",--67
    "0000000000010111",--68
    "0000000000010111",--69
    "0000000000011000",--70
    "0000000000011000",--71
    "0000000000011000",--72
    "0000000000011001",--73
    "0000000000011001",--74
    "0000000000011010",--75
    "0000000000011010",--76
    "0000000000011011",--77
    "0000000000011011",--78
    "0000000000011100",--79
    "0000000000011100",--80
    "0000000000011101",--81
    "0000000000011101",--82
    "0000000000011101",--83
    "0000000000011110",--84
    "0000000000011110",--85
    "0000000000011111",--86
    "0000000000011111",--87
    "0000000000100000",--88
    "0000000000100000",--89
    "0000000000100001",--90
    "0000000000100001",--91
    "0000000000100010",--92
    "0000000000100010",--93
    "0000000000100011",--94
    "0000000000100011",--95
    "0000000000100100",--96
    "0000000000100100",--97
    "0000000000100101",--98
    "0000000000100110",--99
    "0000000000100110",--100
    "0000000000100111",--101
    "0000000000100111",--102
    "0000000000101000",--103
    "0000000000101000",--104
    "0000000000101001",--105
    "0000000000101001",--106
    "0000000000101010",--107
    "0000000000101010",--108
    "0000000000101011",--109
    "0000000000101011",--110
    "0000000000101100",--111
    "0000000000101101",--112
    "0000000000101101",--113
    "0000000000101110",--114
    "0000000000101110",--115
    "0000000000101111",--116
    "0000000000101111",--117
    "0000000000110000",--118
    "0000000000110000",--119
    "0000000000110001",--120
    "0000000000110010",--121
    "0000000000110010",--122
    "0000000000110011",--123
    "0000000000110011",--124
    "0000000000110100",--125
    "0000000000110100",--126
    "0000000000110101",--127
    "0000000000110110",--128
    "0000000000110110",--129
    "0000000000110111",--130
    "0000000000110111",--131
    "0000000000111000",--132
    "0000000000111000",--133
    "0000000000111001",--134
    "0000000000111010",--135
    "0000000000111010",--136
    "0000000000111011",--137
    "0000000000111011",--138
    "0000000000111100",--139
    "0000000000111100",--140
    "0000000000111101",--141
    "0000000000111101",--142
    "0000000000111110",--143
    "0000000000111111",--144
    "0000000000111111",--145
    "0000000001000000",--146
    "0000000001000000",--147
    "0000000001000001",--148
    "0000000001000001",--149
    "0000000001000010",--150
    "0000000001000010",--151
    "0000000001000011",--152
    "0000000001000100",--153
    "0000000001000100",--154
    "0000000001000101",--155
    "0000000001000101",--156
    "0000000001000110",--157
    "0000000001000110",--158
    "0000000001000111",--159
    "0000000001000111",--160
    "0000000001001000",--161
    "0000000001001000",--162
    "0000000001001001",--163
    "0000000001001001",--164
    "0000000001001010",--165
    "0000000001001010",--166
    "0000000001001011",--167
    "0000000001001011",--168
    "0000000001001100",--169
    "0000000001001100",--170
    "0000000001001101",--171
    "0000000001001101",--172
    "0000000001001110",--173
    "0000000001001110",--174
    "0000000001001111",--175
    "0000000001001111",--176
    "0000000001010000",--177
    "0000000001010000",--178
    "0000000001010001",--179
    "0000000001010001",--180
    "0000000001010010",--181
    "0000000001010010",--182
    "0000000001010010",--183
    "0000000001010011",--184
    "0000000001010011",--185
    "0000000001010100",--186
    "0000000001010100",--187
    "0000000001010101",--188
    "0000000001010101",--189
    "0000000001010101",--190
    "0000000001010110",--191
    "0000000001010110",--192
    "0000000001010111",--193
    "0000000001010111",--194
    "0000000001010111",--195
    "0000000001011000",--196
    "0000000001011000",--197
    "0000000001011001",--198
    "0000000001011001",--199
    "0000000001011001",--200
    "0000000001011010",--201
    "0000000001011010",--202
    "0000000001011010",--203
    "0000000001011011",--204
    "0000000001011011",--205
    "0000000001011011",--206
    "0000000001011100",--207
    "0000000001011100",--208
    "0000000001011100",--209
    "0000000001011101",--210
    "0000000001011101",--211
    "0000000001011101",--212
    "0000000001011110",--213
    "0000000001011110",--214
    "0000000001011110",--215
    "0000000001011110",--216
    "0000000001011111",--217
    "0000000001011111",--218
    "0000000001011111",--219
    "0000000001011111",--220
    "0000000001100000",--221
    "0000000001100000",--222
    "0000000001100000",--223
    "0000000001100000",--224
    "0000000001100001",--225
    "0000000001100001",--226
    "0000000001100001",--227
    "0000000001100001",--228
    "0000000001100001",--229
    "0000000001100010",--230
    "0000000001100010",--231
    "0000000001100010",--232
    "0000000001100010",--233
    "0000000001100010",--234
    "0000000001100010",--235
    "0000000001100011",--236
    "0000000001100011",--237
    "0000000001100011",--238
    "0000000001100011",--239
    "0000000001100011",--240
    "0000000001100011",--241
    "0000000001100011",--242
    "0000000001100011",--243
    "0000000001100011",--244
    "0000000001100100",--245
    "0000000001100100",--246
    "0000000001100100",--247
    "0000000001100100",--248
    "0000000001100100",--249
    "0000000001100100",--250
    "0000000001100100",--251
    "0000000001100100",--252
    "0000000001100100",--253
    "0000000001100100",--254
    "0000000001100100",--255
    "0000000001100100",--256
    "0000000001100100",--257
    "0000000001100100",--258
    "0000000001100100",--259
    "0000000001100100",--260
    "0000000001100100",--261
    "0000000001100100",--262
    "0000000001100100",--263
    "0000000001100100",--264
    "0000000001100100",--265
    "0000000001100100",--266
    "0000000001100100",--267
    "0000000001100100",--268
    "0000000001100011",--269
    "0000000001100011",--270
    "0000000001100011",--271
    "0000000001100011",--272
    "0000000001100011",--273
    "0000000001100011",--274
    "0000000001100011",--275
    "0000000001100011",--276
    "0000000001100011",--277
    "0000000001100010",--278
    "0000000001100010",--279
    "0000000001100010",--280
    "0000000001100010",--281
    "0000000001100010",--282
    "0000000001100010",--283
    "0000000001100001",--284
    "0000000001100001",--285
    "0000000001100001",--286
    "0000000001100001",--287
    "0000000001100001",--288
    "0000000001100000",--289
    "0000000001100000",--290
    "0000000001100000",--291
    "0000000001100000",--292
    "0000000001011111",--293
    "0000000001011111",--294
    "0000000001011111",--295
    "0000000001011111",--296
    "0000000001011110",--297
    "0000000001011110",--298
    "0000000001011110",--299
    "0000000001011110",--300
    "0000000001011101",--301
    "0000000001011101",--302
    "0000000001011101",--303
    "0000000001011100",--304
    "0000000001011100",--305
    "0000000001011100",--306
    "0000000001011011",--307
    "0000000001011011",--308
    "0000000001011011",--309
    "0000000001011010",--310
    "0000000001011010",--311
    "0000000001011010",--312
    "0000000001011001",--313
    "0000000001011001",--314
    "0000000001011001",--315
    "0000000001011000",--316
    "0000000001011000",--317
    "0000000001010111",--318
    "0000000001010111",--319
    "0000000001010111",--320
    "0000000001010110",--321
    "0000000001010110",--322
    "0000000001010101",--323
    "0000000001010101",--324
    "0000000001010101",--325
    "0000000001010100",--326
    "0000000001010100",--327
    "0000000001010011",--328
    "0000000001010011",--329
    "0000000001010010",--330
    "0000000001010010",--331
    "0000000001010010",--332
    "0000000001010001",--333
    "0000000001010001",--334
    "0000000001010000",--335
    "0000000001010000",--336
    "0000000001001111",--337
    "0000000001001111",--338
    "0000000001001110",--339
    "0000000001001110",--340
    "0000000001001101",--341
    "0000000001001101",--342
    "0000000001001100",--343
    "0000000001001100",--344
    "0000000001001011",--345
    "0000000001001011",--346
    "0000000001001010",--347
    "0000000001001010",--348
    "0000000001001001",--349
    "0000000001001001",--350
    "0000000001001000",--351
    "0000000001001000",--352
    "0000000001000111",--353
    "0000000001000111",--354
    "0000000001000110",--355
    "0000000001000110",--356
    "0000000001000101",--357
    "0000000001000101",--358
    "0000000001000100",--359
    "0000000001000100",--360
    "0000000001000011",--361
    "0000000001000010",--362
    "0000000001000010",--363
    "0000000001000001",--364
    "0000000001000001",--365
    "0000000001000000",--366
    "0000000001000000",--367
    "0000000000111111",--368
    "0000000000111111",--369
    "0000000000111110",--370
    "0000000000111101",--371
    "0000000000111101",--372
    "0000000000111100",--373
    "0000000000111100",--374
    "0000000000111011",--375
    "0000000000111011",--376
    "0000000000111010",--377
    "0000000000111010",--378
    "0000000000111001",--379
    "0000000000111000",--380
    "0000000000111000",--381
    "0000000000110111",--382
    "0000000000110111",--383
    "0000000000110110",--384
    "0000000000110110",--385
    "0000000000110101",--386
    "0000000000110100",--387
    "0000000000110100",--388
    "0000000000110011",--389
    "0000000000110011",--390
    "0000000000110010",--391
    "0000000000110010",--392
    "0000000000110001",--393
    "0000000000110000",--394
    "0000000000110000",--395
    "0000000000101111",--396
    "0000000000101111",--397
    "0000000000101110",--398
    "0000000000101110",--399
    "0000000000101101",--400
    "0000000000101101",--401
    "0000000000101100",--402
    "0000000000101011",--403
    "0000000000101011",--404
    "0000000000101010",--405
    "0000000000101010",--406
    "0000000000101001",--407
    "0000000000101001",--408
    "0000000000101000",--409
    "0000000000101000",--410
    "0000000000100111",--411
    "0000000000100111",--412
    "0000000000100110",--413
    "0000000000100110",--414
    "0000000000100101",--415
    "0000000000100100",--416
    "0000000000100100",--417
    "0000000000100011",--418
    "0000000000100011",--419
    "0000000000100010",--420
    "0000000000100010",--421
    "0000000000100001",--422
    "0000000000100001",--423
    "0000000000100000",--424
    "0000000000100000",--425
    "0000000000011111",--426
    "0000000000011111",--427
    "0000000000011110",--428
    "0000000000011110",--429
    "0000000000011101",--430
    "0000000000011101",--431
    "0000000000011101",--432
    "0000000000011100",--433
    "0000000000011100",--434
    "0000000000011011",--435
    "0000000000011011",--436
    "0000000000011010",--437
    "0000000000011010",--438
    "0000000000011001",--439
    "0000000000011001",--440
    "0000000000011000",--441
    "0000000000011000",--442
    "0000000000011000",--443
    "0000000000010111",--444
    "0000000000010111",--445
    "0000000000010110",--446
    "0000000000010110",--447
    "0000000000010110",--448
    "0000000000010101",--449
    "0000000000010101",--450
    "0000000000010100",--451
    "0000000000010100",--452
    "0000000000010100",--453
    "0000000000010011",--454
    "0000000000010011",--455
    "0000000000010010",--456
    "0000000000010010",--457
    "0000000000010010",--458
    "0000000000010001",--459
    "0000000000010001",--460
    "0000000000010001",--461
    "0000000000010000",--462
    "0000000000010000",--463
    "0000000000010000",--464
    "0000000000001111",--465
    "0000000000001111",--466
    "0000000000001111",--467
    "0000000000001111",--468
    "0000000000001110",--469
    "0000000000001110",--470
    "0000000000001110",--471
    "0000000000001101",--472
    "0000000000001101",--473
    "0000000000001101",--474
    "0000000000001101",--475
    "0000000000001100",--476
    "0000000000001100",--477
    "0000000000001100",--478
    "0000000000001100",--479
    "0000000000001100",--480
    "0000000000001011",--481
    "0000000000001011",--482
    "0000000000001011",--483
    "0000000000001011",--484
    "0000000000001011",--485
    "0000000000001010",--486
    "0000000000001010",--487
    "0000000000001010",--488
    "0000000000001010",--489
    "0000000000001010",--490
    "0000000000001010",--491
    "0000000000001001",--492
    "0000000000001001",--493
    "0000000000001001",--494
    "0000000000001001",--495
    "0000000000001001",--496
    "0000000000001001",--497
    "0000000000001001",--498
    "0000000000001001",--499
    "0000000000001000",--500
    "0000000000001000",--501
    "0000000000001000",--502
    "0000000000001000",--503
    "0000000000001000",--504
    "0000000000001000",--505
    "0000000000001000",--506
    "0000000000001000",--507
    "0000000000001000",--508
    "0000000000001000",--509
    "0000000000001000",--510
    "0000000000001000",--511
    "0000000000001000");--512


begin

data<=rom(address);

end Behavioral;